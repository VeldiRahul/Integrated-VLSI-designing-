interface vmc_if(input logic clk);
  logic rstn;
  logic cfg_mode;
endinterface

