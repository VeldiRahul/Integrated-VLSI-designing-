interface currency_if(input logic clk);
  logic        currency_valid;
  logic [7:0]  currency_value; 
endinterface